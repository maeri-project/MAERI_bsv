typedef 16 DistributionBandwidth;
typedef 16 CollectionBandwidth;
typedef 128 NumMultSwitches;
